///////////////////////////////////////////////////////
// seg_decoder.v
//
// 기능: 4비트 입력(digit)을 받아 해당하는 숫자/문자를 7세그먼트 형식으로 디코딩
//
// 매핑:
// 0~9 : 숫자 표시
// A, L, I, F, '-' : 문자 표시
// 디코딩 결과를 seg로 출력 (a~g 세그먼트 활성화)
//
// 입력:
// - digit : 표시하고자 하는 값(0~9, A=10, L=11, I=12, F=13, '-'=14)
//
// 출력:
// - seg : 해당 digit에 대응하는 7세그먼트 패턴 (active low 방식)
//
// 참고:
// '1'과 유사한 I, 'L'은 간단히 특정 패턴으로 표시
///////////////////////////////////////////////////////
module seg_decoder(
    input [3:0] digit,
    output reg [6:0] seg
    );
    always @(*) begin
        case(digit)
            4'd0: seg = 7'b1000000; //0
            4'd1: seg = 7'b1111001; //1
            4'd2: seg = 7'b0100100; //2
            4'd3: seg = 7'b0110000; //3
            4'd4: seg = 7'b0011001; //4
            4'd5: seg = 7'b0010010; //5
            4'd6: seg = 7'b0000010; //6
            4'd7: seg = 7'b1111000; //7
            4'd8: seg = 7'b0000000; //8
            4'd9: seg = 7'b0010000; //9
            4'ha: seg = 7'b0001000; //A
            4'hb: seg = 7'b1000111; //L
            4'hc: seg = 7'b1111001; //I (1 형태)
            4'hd: seg = 7'b0001110; //F
            4'he: seg = 7'b0111111; //'-'
            default: seg = 7'b1111111; // default: all off
        endcase
    end
endmodule
